module SubText(
    input               clk,
    input   [95:0]      az, bz, z,
    input   [63:0]      a, b,
    output  [63:0]      aq, bq
    );
    
    wire[63:0] res_a, res_b;
    
    SBox sbox0   (  .clk(clk), .A(a[63:60]), .B(b[63:60]), .A_out(res_a[63:60]), .B_out(res_b[63:60]), 
                    .Az0(az[95:94]), .Az1(az[93:92]), .Az2(az[91:90]), 
                    .Bz0(bz[95:94]), .Bz1(bz[93:92]), .Bz2(bz[91:90]), 
                     .Z0( z[95:94]),  .Z1( z[93:92]),  .Z2( z[91:90]));
                    
    SBox sbox1   (  .clk(clk), .A(a[59:56]), .B(b[59:56]), .A_out(res_a[59:56]), .B_out(res_b[59:56]), 
                    .Az0(az[89:88]), .Az1(az[87:86]), .Az2(az[85:84]), 
                    .Bz0(bz[89:88]), .Bz1(bz[87:86]), .Bz2(bz[85:84]), 
                     .Z0( z[89:88]),  .Z1( z[87:86]),  .Z2( z[85:84]));
                    
    SBox sbox2   (  .clk(clk), .A(a[55:52]), .B(b[55:52]), .A_out(res_a[55:52]), .B_out(res_b[55:52]), 
                    .Az0(az[83:82]), .Az1(az[81:80]), .Az2(az[79:78]), 
                    .Bz0(bz[83:82]), .Bz1(bz[81:80]), .Bz2(bz[79:78]), 
                     .Z0( z[83:82]),  .Z1( z[81:80]),  .Z2( z[79:78]));
                    
    SBox sbox3   (  .clk(clk), .A(a[51:48]), .B(b[51:48]), .A_out(res_a[51:48]), .B_out(res_b[51:48]), 
                    .Az0(az[77:76]), .Az1(az[75:74]), .Az2(az[73:72]), 
                    .Bz0(bz[77:76]), .Bz1(bz[75:74]), .Bz2(bz[73:72]), 
                     .Z0( z[77:76]),  .Z1( z[75:74]),  .Z2( z[73:72]));
                    
    SBox sbox4   (  .clk(clk), .A(a[47:44]), .B(b[47:44]), .A_out(res_a[47:44]), .B_out(res_b[47:44]), 
                    .Az0(az[71:70]), .Az1(az[69:68]), .Az2(az[67:66]), 
                    .Bz0(bz[71:70]), .Bz1(bz[69:68]), .Bz2(bz[67:66]), 
                     .Z0( z[71:70]),  .Z1( z[69:68]),  .Z2( z[67:66]));
                    
    SBox sbox5   (  .clk(clk), .A(a[43:40]), .B(b[43:40]), .A_out(res_a[43:40]), .B_out(res_b[43:40]), 
                    .Az0(az[65:64]), .Az1(az[63:62]), .Az2(az[61:60]), 
                    .Bz0(bz[65:64]), .Bz1(bz[63:62]), .Bz2(bz[61:60]), 
                     .Z0( z[65:64]),  .Z1( z[63:62]),  .Z2( z[61:60]));
                    
    SBox sbox6   (  .clk(clk), .A(a[39:36]), .B(b[39:36]), .A_out(res_a[39:36]), .B_out(res_b[39:36]), 
                    .Az0(az[59:58]), .Az1(az[57:56]), .Az2(az[55:54]), 
                    .Bz0(bz[59:58]), .Bz1(bz[57:56]), .Bz2(bz[55:54]), 
                     .Z0( z[59:58]),  .Z1( z[57:56]),  .Z2( z[55:54]));
                    
    SBox sbox7   (  .clk(clk), .A(a[35:32]), .B(b[35:32]), .A_out(res_a[35:32]), .B_out(res_b[35:32]), 
                    .Az0(az[53:52]), .Az1(az[51:50]), .Az2(az[49:48]), 
                    .Bz0(bz[53:52]), .Bz1(bz[51:50]), .Bz2(bz[49:48]), 
                     .Z0( z[53:52]),  .Z1( z[51:50]),  .Z2( z[49:48])); 
                    
    SBox sbox8   (  .clk(clk), .A(a[31:28]), .B(b[31:28]), .A_out(res_a[31:28]), .B_out(res_b[31:28]), 
                    .Az0(az[47:46]), .Az1(az[45:44]), .Az2(az[43:42]), 
                    .Bz0(bz[47:46]), .Bz1(bz[45:44]), .Bz2(bz[43:42]), 
                     .Z0( z[47:46]),  .Z1( z[45:44]),  .Z2( z[43:42])); 
                    
    SBox sbox9   (  .clk(clk), .A(a[27:24]), .B(b[27:24]), .A_out(res_a[27:24]), .B_out(res_b[27:24]), 
                    .Az0(az[41:40]), .Az1(az[39:38]), .Az2(az[37:36]), 
                    .Bz0(bz[41:40]), .Bz1(bz[39:38]), .Bz2(bz[37:36]), 
                     .Z0( z[41:40]),  .Z1( z[39:38]),  .Z2( z[37:36]));
                    
    SBox sbox10  (  .clk(clk), .A(a[23:20]), .B(b[23:20]), .A_out(res_a[23:20]), .B_out(res_b[23:20]), 
                    .Az0(az[35:34]), .Az1(az[33:32]), .Az2(az[31:30]), 
                    .Bz0(bz[35:34]), .Bz1(bz[33:32]), .Bz2(bz[31:30]), 
                     .Z0( z[35:34]),  .Z1( z[33:32]),  .Z2( z[31:30]));
                    
    SBox sbox11  (  .clk(clk), .A(a[19:16]), .B(b[19:16]), .A_out(res_a[19:16]), .B_out(res_b[19:16]), 
                    .Az0(az[29:28]), .Az1(az[27:26]), .Az2(az[25:24]), 
                    .Bz0(bz[29:28]), .Bz1(bz[27:26]), .Bz2(bz[25:24]), 
                     .Z0( z[29:28]),  .Z1( z[27:26]),  .Z2( z[25:24]));
                    
    SBox sbox12  (  .clk(clk), .A(a[15:12]), .B(b[15:12]), .A_out(res_a[15:12]), .B_out(res_b[15:12]), 
                    .Az0(az[23:22]), .Az1(az[21:20]), .Az2(az[19:18]), 
                    .Bz0(bz[23:22]), .Bz1(bz[21:20]), .Bz2(bz[19:18]), 
                     .Z0( z[23:22]),  .Z1( z[21:20]),  .Z2( z[19:18]));
                    
    SBox sbox13  (  .clk(clk), .A(a[11:08]), .B(b[11:08]), .A_out(res_a[11:08]), .B_out(res_b[11:08]), 
                    .Az0(az[17:16]), .Az1(az[15:14]), .Az2(az[13:12]), 
                    .Bz0(bz[17:16]), .Bz1(bz[15:14]), .Bz2(bz[13:12]), 
                     .Z0( z[17:16]),  .Z1( z[15:14]),  .Z2( z[13:12]));
                    
    SBox sbox14  (  .clk(clk), .A(a[07:04]), .B(b[07:04]), .A_out(res_a[07:04]), .B_out(res_b[07:04]), 
                    .Az0(az[11:10]), .Az1(az[09:08]), .Az2(az[07:06]), 
                    .Bz0(bz[11:10]), .Bz1(bz[09:08]), .Bz2(bz[07:06]), 
                     .Z0( z[11:10]),  .Z1( z[09:08]),  .Z2( z[07:06]));
                    
    SBox sbox15  (  .clk(clk), .A(a[03:00]), .B(b[03:00]), .A_out(res_a[03:00]), .B_out(res_b[03:00]), 
                    .Az0(az[05:04]), .Az1(az[03:02]), .Az2(az[01:00]), 
                    .Bz0(bz[05:04]), .Bz1(bz[03:02]), .Bz2(bz[01:00]), 
                     .Z0( z[05:04]),  .Z1( z[03:02]),  .Z2( z[01:00])); 
                    
    assign aq = res_a;
    assign bq = res_b;
                   
endmodule